module not_gate(
    input A_i,
    output F_o
);
    assign F_o = ~A_i;
endmodule